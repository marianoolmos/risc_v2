--====================================================================
--
--   /@@@@@@@  /@@@@@@  /@@@@@@   /@@@@@@        /@@    /@@  /@@@@@@
--  | @@__  @@|_  @@_/ /@@__  @@ /@@__  @@      | @@   | @@ /@@__  @@
--  | @@  \ @@  | @@  | @@  \__/| @@  \__/      | @@   | @@|__/  \ @@
--  | @@@@@@@/  | @@  |  @@@@@@ | @@            |  @@ / @@/  /@@@@@@/
--  | @@__  @@  | @@   \____  @@| @@             \  @@ @@/  /@@____/
--  | @@  \ @@  | @@   /@@  \ @@| @@    @@        \  @@@/  | @@
--  | @@  | @@ /@@@@@@|  @@@@@@/|  @@@@@@/         \  @/   | @@@@@@@@
--  |__/  |__/|______/ \______/  \______/           \_/    |________/
--
-- Module:       RISC_V2_REG_FILE
-- Description:
--
-- Author:       Mariano Olmos Martin
-- Mail  :       mariano.olmos@outlook.com
-- Date:         13/9/2025
-- Version:      v0.0
-- License: MIT License
--
-- Copyright (c) 2025 Mariano Olmos
--
-- Permission is hereby granted, free of charge, to any person obtaining
-- a copy of this VHDL code and associated documentation files (the
-- "Software"), to deal in the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject
-- to the following conditions:
--
-- The above copyright notice and this permission notice shall be
-- included in all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
-- OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
-- NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS BE LIABLE FOR ANY
-- CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
--======================================================================

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
  use ieee.math_real.all;
  use work.risc_v2_pkg.all;

entity risc_v2_reg_file is
  port (
    clk   : in    std_logic;
    reset : in    std_logic;
    we    : in    std_logic;
    rs1   : in    std_logic_vector(31 downto 0);
    rs2   : in    std_logic_vector(31 downto 0);
    din   : in    std_logic_vector(31 downto 0);
    rd    : in    std_logic_vector(31 downto 0);
    dout1 : out   std_logic_vector(31 downto 0);
    dout2 : out   std_logic_vector(31 downto 0)
  );
end entity risc_v2_reg_file;

architecture rtl of risc_v2_reg_file is

  type rf_t is array(0 to 2 ** rd'length - 1) of std_logic_vector(din'length - 1 downto 0);

  signal rf : rf_t;

begin

  process (clk, reset) is
  begin

    if (reset = '1') then
      rf <= (others => (others => '0'));
    elsif rising_edge(clk) then
      if (we = '1') then
        rf(to_integer(unsigned(rd))) <= din;
      end if;
    end if;

  end process;

  -- Escritura síncrona
  dout1 <= rf(to_integer(unsigned(rs1))); -- Lectura asíncrona
  dout2 <= rf(to_integer(unsigned(rs2))); -- Lectura asíncrona

end architecture rtl;
